`timescale 1 ns / 1 ps
`include "alu.v"

module testALU();
    
    reg[31:0] a;
    reg[31:0] b;

    wire[31:0] out;
    wire overflow;

endmodule

