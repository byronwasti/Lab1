// define logic control
`define ADD  3'd0
`define SUB  3'd1
`define XOR  3'd2
`define SLT  3'd3
`define AND  3'd4
`define NAND 3'd5
`define NOR  3'd6
`define OR   3'd7


module aluLUT
(
    output reg[2:0] sel,
    output reg      negate,
    input[2:0]      ALUcommand
)

  always// @(ALUcommand) 
  begin
    case (ALUcommand)
        `ADD:  begin muxindex = 0; invert=0; end    
        `SUB:  begin muxindex = 0; invert=1; end
        `AND:  begin muxindex = 1; invert=1; end
        `NAND: begin muxindex = 1; invert=0; end
        `NOR:  begin muxindex = 2; invert=0; end
        `OR:   begin muxindex = 2; invert=1; end
        `XOR:  begin muxindex = 3; invert=0; end
        // `SLT:  begin muxindex = 2; invert=0; end   
    endcase
  end
endmodule
